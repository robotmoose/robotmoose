** Profile: "SCHEMATIC1-AC Sweep"  [ C:\Users\Ryker Dial\Documents\Documents\UAF\Robotics\ITEST\Sound Localization Research\OrCAD\wide_bandpass-pspicefiles\schematic1\ac sweep.sim ] 

** Creating circuit file "AC Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Ryker Dial\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 
.lib "fairchild.lib" 
.lib "bipolar.lib" 
.lib "diode.lib" 

*Analysis directives: 
.AC DEC 100 10 100k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

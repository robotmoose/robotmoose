** Profile: "SCHEMATIC1-wfea"  [ C:\OrCAD_Projects\Wide_BandPass-PSpiceFiles\SCHEMATIC1\wfea.sim ] 

** Creating circuit file "wfea.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Ryker Dial\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 
.lib "fairchild.lib" 
.lib "bipolar.lib" 
.lib "diode.lib" 

*Analysis directives: 
.AC DEC 100 100m 100k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
